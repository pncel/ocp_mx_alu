
module mx_alu (
    // TODO top-level interface of the whole ALU
);

    // TODO parsing top-level interface into appropriate functional units

endmodule