
`ifndef ALU_CORE_PKG
`define ALU_CORE_PKG

package alu_core_pkg;
    import alu_op_pkg::*;
    import mx_format_pkg::*;
    import mx_function_pkg::*;
    import scalar_format_pkg::*;
endpackage

`endif // ALU_CORE_PKG